library verilog;
use verilog.vl_types.all;
entity MUX_2_1_8BITS_vlg_vec_tst is
end MUX_2_1_8BITS_vlg_vec_tst;
