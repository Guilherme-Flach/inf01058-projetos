library verilog;
use verilog.vl_types.all;
entity ULA4bits_vlg_vec_tst is
end ULA4bits_vlg_vec_tst;
