library verilog;
use verilog.vl_types.all;
entity FREQ_DIV_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FREQ_DIV_vlg_check_tst;
