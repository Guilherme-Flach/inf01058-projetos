library verilog;
use verilog.vl_types.all;
entity DEC_16_vlg_vec_tst is
end DEC_16_vlg_vec_tst;
