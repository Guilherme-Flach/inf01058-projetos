library verilog;
use verilog.vl_types.all;
entity FREQ_DIV_vlg_vec_tst is
end FREQ_DIV_vlg_vec_tst;
