library verilog;
use verilog.vl_types.all;
entity LAB01_vlg_vec_tst is
end LAB01_vlg_vec_tst;
