library verilog;
use verilog.vl_types.all;
entity PROJETO_NEANDER_RAM_vlg_vec_tst is
end PROJETO_NEANDER_RAM_vlg_vec_tst;
