library verilog;
use verilog.vl_types.all;
entity PROJETO_NEANDER_RAM_vlg_check_tst is
    port(
        AC0_A           : in     vl_logic;
        AC0_B           : in     vl_logic;
        AC0_C           : in     vl_logic;
        AC0_D           : in     vl_logic;
        AC0_E           : in     vl_logic;
        AC0_F           : in     vl_logic;
        AC0_G           : in     vl_logic;
        AC1_A           : in     vl_logic;
        AC1_B           : in     vl_logic;
        AC1_C           : in     vl_logic;
        AC1_D           : in     vl_logic;
        AC1_E           : in     vl_logic;
        AC1_F           : in     vl_logic;
        AC1_G           : in     vl_logic;
        AC_O            : in     vl_logic_vector(7 downto 0);
        ADDR            : in     vl_logic_vector(7 downto 0);
        C_AC            : in     vl_logic;
        C_NZ            : in     vl_logic;
        C_PC            : in     vl_logic;
        C_RDM           : in     vl_logic;
        C_REM           : in     vl_logic;
        C_RI            : in     vl_logic;
        DATA            : in     vl_logic_vector(7 downto 0);
        GOTO_T0         : in     vl_logic;
        HLT_OUT         : in     vl_logic;
        INC_PC          : in     vl_logic;
        N_OUT           : in     vl_logic;
        PC0_A           : in     vl_logic;
        PC0_B           : in     vl_logic;
        PC0_C           : in     vl_logic;
        PC0_D           : in     vl_logic;
        PC0_E           : in     vl_logic;
        PC0_F           : in     vl_logic;
        PC0_G           : in     vl_logic;
        PC1_A           : in     vl_logic;
        PC1_B           : in     vl_logic;
        PC1_C           : in     vl_logic;
        PC1_D           : in     vl_logic;
        PC1_E           : in     vl_logic;
        PC1_F           : in     vl_logic;
        PC1_G           : in     vl_logic;
        PC_O            : in     vl_logic_vector(7 downto 0);
        READ            : in     vl_logic;
        RI_O            : in     vl_logic_vector(7 downto 0);
        SEL             : in     vl_logic;
        TEMP_O          : in     vl_logic_vector(7 downto 0);
        ULA_ADD         : in     vl_logic;
        ULA_AND         : in     vl_logic;
        ULA_NOT         : in     vl_logic;
        ULA_OR          : in     vl_logic;
        ULA_Y           : in     vl_logic;
        WRITE           : in     vl_logic;
        Z_OUT           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end PROJETO_NEANDER_RAM_vlg_check_tst;
