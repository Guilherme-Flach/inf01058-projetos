library verilog;
use verilog.vl_types.all;
entity CONT_UP_DOWN_vlg_vec_tst is
end CONT_UP_DOWN_vlg_vec_tst;
