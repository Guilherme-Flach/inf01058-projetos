library verilog;
use verilog.vl_types.all;
entity CONT_UP_DOWN_vlg_check_tst is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        E0              : in     vl_logic;
        E1              : in     vl_logic;
        F0              : in     vl_logic;
        F1              : in     vl_logic;
        G0              : in     vl_logic;
        G1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CONT_UP_DOWN_vlg_check_tst;
